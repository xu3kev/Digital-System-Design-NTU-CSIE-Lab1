module full_adder(a, b, sum, cin, cout);

input a;
input b;
input cin;
output sum;
output cout;
/*
TODO:
use gate level primitives to construct a full adder
Useful gate primitives: or, and , xor
*/

endmodule
