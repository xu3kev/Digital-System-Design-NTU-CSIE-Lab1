module binary_adder( a, b, sum);
input [5:0] a;
input [5:0] b;
output [5:0] sum;
/*
TODO:
use full_adder module to build a binary adder:
a + b = sum
Please see the testbench binary_adder_tb.v for the sample input and output.
*/

endmodule
